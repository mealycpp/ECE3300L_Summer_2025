module decoder4x16_gate (

);
endmodule