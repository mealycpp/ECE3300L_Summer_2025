module tb_decoder4x16 (

);
endmodule