module decoder4x16_Behavior (
  input  wire [3:0] I,
    input  wire       W,
  output reg  [15:0] O
);

always @(*) begin
  //reseting to 0
    O = 16'b0; 
  // only decoding if enabled is the catch
  if (W) begin 
    case (I)
            4'b0000: O = 16'b0000_0000_0000_0001; 
            4'b0001: O = 16'b0000_0000_0000_0010;
            4'b0010: O = 16'b0000_0000_0000_0100;
            4'b0011: O = 16'b0000_0000_0000_1000;
            4'b0100: O = 16'b0000_0000_0001_0000;
            4'b0101: O = 16'b0000_0000_0010_0000;
            4'b0110: O = 16'b0000_0000_0100_0000;
            4'b0111: O = 16'b0000_0000_1000_0000;
            4'b1000: O = 16'b0000_0001_0000_0000;
            4'b1001: O = 16'b0000_0010_0000_0000;
            4'b1010: O = 16'b0000_0100_0000_0000;
            4'b1011: O = 16'b0000_1000_0000_0000;
            4'b1100: O = 16'b0001_0000_0000_0000;
            4'b1101: O = 16'b0010_0000_0000_0000;
            4'b1110: O = 16'b0100_0000_0000_0000;
            4'b1111: O = 16'b1000_0000_0000_0000;
        endcase
    end
end

endmodule
