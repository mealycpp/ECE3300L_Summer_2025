`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/11/2025 01:09:04 AM
// Design Name: 
// Module Name: ECE3300Lproject1_code
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ECE3300Lproject1_code(
input wire [15:0] sw,
output wire [15:0] led
);
assign led = sw;
endmodule

