`timescale 1ns/1ps
module clock_divider_fixed #(
    parameter integer INPUT_HZ = 100_000_000,
    parameter integer TICK1_HZ = 1_000,
    parameter integer PWM_HZ   = 20_000
)(
    input wire clk_in,
    input wire rst_n,
    output reg clk_1k,
    output reg clk_pwm
);

localparam integer DIV1H  = (INPUT_HZ / TICK1_HZ) / 2;
localparam integer DIVPMH = (INPUT_HZ / PWM_HZ) / 2;

localparam integer WIDTH1  = $clog2(DIV1H);
localparam integer WIDTHPM = $clog2(DIVPMH);

reg [WIDTH1-1:0]  c1;
reg [WIDTHPM-1:0] c2;

always @(posedge clk_in or negedge rst_n) begin
    if (!rst_n) begin
        c1       <= 0;
        clk_1k   <= 0;
        c2       <= 0;
        clk_pwm  <= 0;
    end else begin
        // 1 kHz clock toggle
        if (c1 == DIV1H - 1) begin
            c1     <= 0;
            clk_1k <= ~clk_1k;
        end else begin
            c1 <= c1 + 1;
        end

        // 20 kHz clock toggle
        if (c2 == DIVPMH - 1) begin
            c2      <= 0;
            clk_pwm <= ~clk_pwm;
        end else begin
            c2 <= c2 + 1;
        end
    end
end

endmodule
