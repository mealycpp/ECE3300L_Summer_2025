module decoder4x16_behav (
    input [4:0] sw,
    output reg [15:0] led
);
    always @(*) begin
        led = 16'b0; // Green Resets outputs to 0
        if (sw[4]) begin // Blue cEheck if enabled
            case (sw[3:0])
                4'b0000: led = 16'b0000_0000_0000_0001; // Output 0
                4'b0001: led = 16'b0000_0000_0000_0010; // Output 1
                4'b0010: led = 16'b0000_0000_0000_0100;
                4'b0011: led = 16'b0000_0000_0000_1000;
                4'b0100: led = 16'b0000_0000_0001_0000;
                4'b0101: led = 16'b0000_0000_0010_0000;
                4'b0110: led = 16'b0000_0000_0100_0000;
                4'b0111: led = 16'b0000_0000_1000_0000;
                4'b1000: led = 16'b0000_0001_0000_0000;
                4'b1001: led = 16'b0000_0010_0000_0000;
                4'b1010: led = 16'b0000_0100_0000_0000;
                4'b1011: led = 16'b0000_1000_0000_0000;
                4'b1100: led = 16'b0001_0000_0000_0000;
                4'b1101: led = 16'b0010_0000_0000_0000;
                4'b1110: led = 16'b0100_0000_0000_0000;
                4'b1111: led = 16'b1000_0000_0000_0000;
            endcase
        end
    end
endmodule