module decoder4x16_behav (

);
endmodule
